module top_module (
    input clk,
    input d, 
    input r,   // synchronous reset
    output q);

endmodule
